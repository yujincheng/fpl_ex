ddr3_nc[0],
ddr3_dq[63],
ddr3_dq[62],
ddr3_dq[61],
ddr3_dq[60],
ddr3_dqs_n[7],
ddr3_dqs_p[7],
ddr3_dq[59],
ddr3_dq[58],
ddr3_dq[57],
ddr3_dq[56],
ddr3_nc[1],
ddr3_dm[7],
ddr3_nc[2],
ddr3_dq[55],
ddr3_dq[54],
ddr3_dq[53],
ddr3_dq[52],
ddr3_dqs_n[6],
ddr3_dqs_p[6],
ddr3_dq[51],
ddr3_dq[50],
ddr3_dq[49],
ddr3_dq[48],
ddr3_nc[3],
ddr3_dm[6],
ddr3_nc[4],
ddr3_dq[47],
ddr3_dq[46],
ddr3_dq[45],
ddr3_dq[44],
ddr3_dqs_n[5],
ddr3_dqs_p[5],
ddr3_dq[43],
ddr3_dq[42],
ddr3_dq[41],
ddr3_dq[40],
ddr3_nc[5],
ddr3_dm[5],
ddr3_nc[6],
ddr3_dq[39],
ddr3_dq[38],
ddr3_dq[37],
ddr3_dq[36],
ddr3_dqs_n[4],
ddr3_dqs_p[4],
ddr3_dq[35],
ddr3_dq[34],
ddr3_dq[33],
ddr3_dq[32],
ddr3_nc[7],
ddr3_dm[4],
ddr3_nc[8],
ddr3_dq[31],
ddr3_dq[30],
ddr3_dq[29],
ddr3_dq[28],
ddr3_dqs_n[3],
ddr3_dqs_p[3],
ddr3_dq[27],
ddr3_dq[26],
ddr3_dq[25],
ddr3_dq[24],
ddr3_nc[9],
ddr3_dm[3],
ddr3_nc[10],
ddr3_dq[23],
ddr3_dq[22],
ddr3_dq[21],
ddr3_dq[20],
ddr3_dqs_n[2],
ddr3_dqs_p[2],
ddr3_dq[19],
ddr3_dq[18],
ddr3_dq[17],
ddr3_dq[16],
ddr3_nc[11],
ddr3_dm[2],
ddr3_nc[12],
ddr3_dq[15],
ddr3_dq[14],
ddr3_dq[13],
ddr3_dq[12],
ddr3_dqs_n[1],
ddr3_dqs_p[1],
ddr3_dq[11],
ddr3_dq[10],
ddr3_dq[9],
ddr3_dq[8],
ddr3_nc[13],
ddr3_dm[1],
ddr3_nc[14],
ddr3_dq[7],
ddr3_dq[6],
ddr3_dq[5],
ddr3_dq[4],
ddr3_dqs_n[0],
ddr3_dqs_p[0],
ddr3_dq[3],
ddr3_dq[2],
ddr3_dq[1],
ddr3_dq[0],
ddr3_nc[15],
ddr3_dm[0],
ddr3_nc[16],
ddr3_nc[17],
ddr3_nc[18],
ddr3_nc[19],
ddr3_nc[20],
ddr3_nc[21],
ddr3_nc[22],
ddr3_nc[23],
ddr3_we_n,
ddr3_cas_n,
ddr3_ras_n,
ddr3_nc[24],
ddr3_odt[0],
ddr3_cke[0],
ddr3_cs_n[0],
ddr3_ba[2],
ddr3_nc[25],
ddr3_nc[26],
ddr3_ba[1],
ddr3_ba[0],
ddr3_addr[15],
ddr3_addr[14],
ddr3_addr[13],
ddr3_addr[12],
ddr3_addr[11],
ddr3_addr[10],
ddr3_nc[27],
ddr3_addr[9],
ddr3_addr[8],
ddr3_addr[7],
ddr3_addr[6],
ddr3_ck_n[0],
ddr3_ck_p[0],
ddr3_addr[5],
ddr3_addr[4],
ddr3_addr[3],
ddr3_addr[2],
ddr3_addr[1],
ddr3_addr[0]
