task init_braminst();
begin
    $readmemh ( "..//sim_data//BP_data//bram_0_0.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[0].BUF_UNIT_2[0].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_0_1.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[0].BUF_UNIT_2[1].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_0_2.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[0].BUF_UNIT_2[2].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_0_3.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[0].BUF_UNIT_2[3].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_1_0.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[1].BUF_UNIT_2[0].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_1_1.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[1].BUF_UNIT_2[1].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_1_2.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[1].BUF_UNIT_2[2].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_1_3.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[1].BUF_UNIT_2[3].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_2_0.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[2].BUF_UNIT_2[0].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_2_1.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[2].BUF_UNIT_2[1].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_2_2.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[2].BUF_UNIT_2[2].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_2_3.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[2].BUF_UNIT_2[3].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_3_0.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[3].BUF_UNIT_2[0].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_3_1.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[3].BUF_UNIT_2[1].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_3_2.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[3].BUF_UNIT_2[2].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_3_3.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[3].BUF_UNIT_2[3].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_4_0.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[4].BUF_UNIT_2[0].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_4_1.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[4].BUF_UNIT_2[1].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_4_2.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[4].BUF_UNIT_2[2].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_4_3.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[4].BUF_UNIT_2[3].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_5_0.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[5].BUF_UNIT_2[0].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_5_1.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[5].BUF_UNIT_2[1].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_5_2.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[5].BUF_UNIT_2[2].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_5_3.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[5].BUF_UNIT_2[3].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_6_0.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[6].BUF_UNIT_2[0].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_6_1.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[6].BUF_UNIT_2[1].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_6_2.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[6].BUF_UNIT_2[2].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_6_3.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[6].BUF_UNIT_2[3].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_7_0.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[7].BUF_UNIT_2[0].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_7_1.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[7].BUF_UNIT_2[1].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_7_2.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[7].BUF_UNIT_2[2].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_7_3.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[7].BUF_UNIT_2[3].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_8_0.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[8].BUF_UNIT_2[0].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_8_1.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[8].BUF_UNIT_2[1].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_8_2.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[8].BUF_UNIT_2[2].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_8_3.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[8].BUF_UNIT_2[3].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_9_0.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[9].BUF_UNIT_2[0].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_9_1.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[9].BUF_UNIT_2[1].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_9_2.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[9].BUF_UNIT_2[2].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_9_3.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[9].BUF_UNIT_2[3].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_10_0.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[10].BUF_UNIT_2[0].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_10_1.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[10].BUF_UNIT_2[1].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_10_2.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[10].BUF_UNIT_2[2].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_10_3.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[10].BUF_UNIT_2[3].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_11_0.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[11].BUF_UNIT_2[0].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_11_1.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[11].BUF_UNIT_2[1].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_11_2.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[11].BUF_UNIT_2[2].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_11_3.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[11].BUF_UNIT_2[3].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_12_0.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[12].BUF_UNIT_2[0].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_12_1.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[12].BUF_UNIT_2[1].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_12_2.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[12].BUF_UNIT_2[2].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_12_3.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[12].BUF_UNIT_2[3].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_13_0.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[13].BUF_UNIT_2[0].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_13_1.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[13].BUF_UNIT_2[1].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_13_2.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[13].BUF_UNIT_2[2].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_13_3.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[13].BUF_UNIT_2[3].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_14_0.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[14].BUF_UNIT_2[0].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_14_1.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[14].BUF_UNIT_2[1].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_14_2.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[14].BUF_UNIT_2[2].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_14_3.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[14].BUF_UNIT_2[3].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_15_0.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[15].BUF_UNIT_2[0].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_15_1.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[15].BUF_UNIT_2[1].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_15_2.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[15].BUF_UNIT_2[2].bram_inst.ram_name);
    $readmemh ( "..//sim_data//BP_data//bram_15_3.txt", sim_tb_top.u_ip_top.cnntop.bp.BUF_UNIT_1[15].BUF_UNIT_2[3].bram_inst.ram_name);
end
endtask
