localparam [MUXCONTROL - 1:0] ST_PAD_INIT_1 = 	 0;
localparam [MUXCONTROL - 1:0] ST_PAD_INIT_2 = 	 1;
localparam [MUXCONTROL - 1:0] ST_PAD_UINIT_1 =  2;
localparam [MUXCONTROL - 1:0] ST_PAD_UINIT_2 =  3;
localparam [MUXCONTROL - 1:0] ST_UPAD_INIT_1 =  4;
localparam [MUXCONTROL - 1:0] ST_UPAD_INIT_2 =  5;
localparam [MUXCONTROL - 1:0] ST_UPAD_UINIT_1 = 6;
localparam [MUXCONTROL - 1:0] ST_UPAD_UINIT_2 = 7;
localparam [MUXCONTROL - 1:0] ST_PAD_INIT_END_1 = 	 8;
localparam [MUXCONTROL - 1:0] ST_PAD_INIT_END_2 = 	 9;
localparam [MUXCONTROL - 1:0] ST_PAD_UINIT_END_1 =  10;
localparam [MUXCONTROL - 1:0] ST_PAD_UINIT_END_2 =  11;
localparam [MUXCONTROL - 1:0] ST_UPAD_INIT_END_1 =  12;
localparam [MUXCONTROL - 1:0] ST_UPAD_INIT_END_2 =  13;
localparam [MUXCONTROL - 1:0] ST_UPAD_UINIT_END_1 = 14;
localparam [MUXCONTROL - 1:0] ST_UPAD_UINIT_END_2 = 15;